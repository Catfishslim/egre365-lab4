entity ALU_TestBench is
end ALU_TestBench;

architecture behavior of ALU_TestBench is

	constant MAX_DELAY : time := 20 ns;
	
	